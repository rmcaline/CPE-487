---will upload file soon
